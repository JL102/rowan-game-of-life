library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VGA is
    port(
        CLOCK_25    :   in std_logic
        
    );

end VGA

architecture rtl